module decoder6to64(encoded, decoded);
	input [5:0] encoded;
	output reg [63:0] decoded;

	always @(*)
	case(encoded)
	6'd0   : decoded = 64'b1 << 1'd0;
	6'd1   : decoded = 64'b1 << 1'd1;
	6'd2   : decoded = 64'b1 << 2'd2;
	6'd3   : decoded = 64'b1 << 2'd3;
	6'd4   : decoded = 64'b1 << 3'd4;
	6'd5   : decoded = 64'b1 << 3'd5;
	6'd6   : decoded = 64'b1 << 3'd6;
	6'd7   : decoded = 64'b1 << 3'd7;
	6'd8   : decoded = 64'b1 << 4'd8;
	6'd9   : decoded = 64'b1 << 4'd9;
	6'd10  : decoded = 64'b1 << 4'd10;
	6'd11  : decoded = 64'b1 << 4'd11;
	6'd12  : decoded = 64'b1 << 4'd12;
	6'd13  : decoded = 64'b1 << 4'd13;
	6'd14  : decoded = 64'b1 << 4'd14;
	6'd15  : decoded = 64'b1 << 4'd15;
	6'd16  : decoded = 64'b1 << 5'd16;
	6'd17  : decoded = 64'b1 << 5'd17;
	6'd18  : decoded = 64'b1 << 5'd18;
	6'd19  : decoded = 64'b1 << 5'd19;
	6'd20  : decoded = 64'b1 << 5'd20;
	6'd21  : decoded = 64'b1 << 5'd21;
	6'd22  : decoded = 64'b1 << 5'd22;
	6'd23  : decoded = 64'b1 << 5'd23;
	6'd24  : decoded = 64'b1 << 5'd24;
	6'd25  : decoded = 64'b1 << 5'd25;
	6'd26  : decoded = 64'b1 << 5'd26;
	6'd27  : decoded = 64'b1 << 5'd27;
	6'd28  : decoded = 64'b1 << 5'd28;
	6'd29  : decoded = 64'b1 << 5'd29;
	6'd30  : decoded = 64'b1 << 5'd30;
	6'd31  : decoded = 64'b1 << 5'd31;
	6'd32  : decoded = 64'b1 << 6'd32;
	6'd33  : decoded = 64'b1 << 6'd33;
	6'd34  : decoded = 64'b1 << 6'd34;
	6'd35  : decoded = 64'b1 << 6'd35;
	6'd36  : decoded = 64'b1 << 6'd36;
	6'd37  : decoded = 64'b1 << 6'd37;
	6'd38  : decoded = 64'b1 << 6'd38;
	6'd39  : decoded = 64'b1 << 6'd39;
	6'd40  : decoded = 64'b1 << 6'd40;
	6'd41  : decoded = 64'b1 << 6'd41;
	6'd42  : decoded = 64'b1 << 6'd42;
	6'd43  : decoded = 64'b1 << 6'd43;
	6'd44  : decoded = 64'b1 << 6'd44;
	6'd45  : decoded = 64'b1 << 6'd45;
	6'd46  : decoded = 64'b1 << 6'd46;
	6'd47  : decoded = 64'b1 << 6'd47;
	6'd48  : decoded = 64'b1 << 6'd48;
	6'd49  : decoded = 64'b1 << 6'd49;
	6'd50  : decoded = 64'b1 << 6'd50;
	6'd51  : decoded = 64'b1 << 6'd51;
	6'd52  : decoded = 64'b1 << 6'd52;
	6'd53  : decoded = 64'b1 << 6'd53;
	6'd54  : decoded = 64'b1 << 6'd54;
	6'd55  : decoded = 64'b1 << 6'd55;
	6'd56  : decoded = 64'b1 << 6'd56;
	6'd57  : decoded = 64'b1 << 6'd57;
	6'd58  : decoded = 64'b1 << 6'd58;
	6'd59  : decoded = 64'b1 << 6'd59;
	6'd60  : decoded = 64'b1 << 6'd60;
	6'd61  : decoded = 64'b1 << 6'd61;
	6'd62  : decoded = 64'b1 << 6'd62;
	6'd63  : decoded = 64'b1 << 6'd63;
	endcase
endmodule
