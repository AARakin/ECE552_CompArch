module decoder7to128(encoded, decoded);
	input [6:0] encoded;
	output reg [127:0] decoded;

	always @(*)
	case(encoded)
	7'd0   : decoded = 128'b1 << 1'd0;
	7'd1   : decoded = 128'b1 << 1'd1;
	7'd2   : decoded = 128'b1 << 2'd2;
	7'd3   : decoded = 128'b1 << 2'd3;
	7'd4   : decoded = 128'b1 << 3'd4;
	7'd5   : decoded = 128'b1 << 3'd5;
	7'd6   : decoded = 128'b1 << 3'd6;
	7'd7   : decoded = 128'b1 << 3'd7;
	7'd8   : decoded = 128'b1 << 4'd8;
	7'd9   : decoded = 128'b1 << 4'd9;
	7'd10  : decoded = 128'b1 << 4'd10;
	7'd11  : decoded = 128'b1 << 4'd11;
	7'd12  : decoded = 128'b1 << 4'd12;
	7'd13  : decoded = 128'b1 << 4'd13;
	7'd14  : decoded = 128'b1 << 4'd14;
	7'd15  : decoded = 128'b1 << 4'd15;
	7'd16  : decoded = 128'b1 << 5'd16;
	7'd17  : decoded = 128'b1 << 5'd17;
	7'd18  : decoded = 128'b1 << 5'd18;
	7'd19  : decoded = 128'b1 << 5'd19;
	7'd20  : decoded = 128'b1 << 5'd20;
	7'd21  : decoded = 128'b1 << 5'd21;
	7'd22  : decoded = 128'b1 << 5'd22;
	7'd23  : decoded = 128'b1 << 5'd23;
	7'd24  : decoded = 128'b1 << 5'd24;
	7'd25  : decoded = 128'b1 << 5'd25;
	7'd26  : decoded = 128'b1 << 5'd26;
	7'd27  : decoded = 128'b1 << 5'd27;
	7'd28  : decoded = 128'b1 << 5'd28;
	7'd29  : decoded = 128'b1 << 5'd29;
	7'd30  : decoded = 128'b1 << 5'd30;
	7'd31  : decoded = 128'b1 << 5'd31;
	7'd32  : decoded = 128'b1 << 6'd32;
	7'd33  : decoded = 128'b1 << 6'd33;
	7'd34  : decoded = 128'b1 << 6'd34;
	7'd35  : decoded = 128'b1 << 6'd35;
	7'd36  : decoded = 128'b1 << 6'd36;
	7'd37  : decoded = 128'b1 << 6'd37;
	7'd38  : decoded = 128'b1 << 6'd38;
	7'd39  : decoded = 128'b1 << 6'd39;
	7'd40  : decoded = 128'b1 << 6'd40;
	7'd41  : decoded = 128'b1 << 6'd41;
	7'd42  : decoded = 128'b1 << 6'd42;
	7'd43  : decoded = 128'b1 << 6'd43;
	7'd44  : decoded = 128'b1 << 6'd44;
	7'd45  : decoded = 128'b1 << 6'd45;
	7'd46  : decoded = 128'b1 << 6'd46;
	7'd47  : decoded = 128'b1 << 6'd47;
	7'd48  : decoded = 128'b1 << 6'd48;
	7'd49  : decoded = 128'b1 << 6'd49;
	7'd50  : decoded = 128'b1 << 6'd50;
	7'd51  : decoded = 128'b1 << 6'd51;
	7'd52  : decoded = 128'b1 << 6'd52;
	7'd53  : decoded = 128'b1 << 6'd53;
	7'd54  : decoded = 128'b1 << 6'd54;
	7'd55  : decoded = 128'b1 << 6'd55;
	7'd56  : decoded = 128'b1 << 6'd56;
	7'd57  : decoded = 128'b1 << 6'd57;
	7'd58  : decoded = 128'b1 << 6'd58;
	7'd59  : decoded = 128'b1 << 6'd59;
	7'd60  : decoded = 128'b1 << 6'd60;
	7'd61  : decoded = 128'b1 << 6'd61;
	7'd62  : decoded = 128'b1 << 6'd62;
	7'd63  : decoded = 128'b1 << 6'd63;
	7'd64  : decoded = 128'b1 << 7'd64;
	7'd65  : decoded = 128'b1 << 7'd65;
	7'd66  : decoded = 128'b1 << 7'd66;
	7'd67  : decoded = 128'b1 << 7'd67;
	7'd68  : decoded = 128'b1 << 7'd68;
	7'd69  : decoded = 128'b1 << 7'd69;
	7'd70  : decoded = 128'b1 << 7'd70;
	7'd71  : decoded = 128'b1 << 7'd71;
	7'd72  : decoded = 128'b1 << 7'd72;
	7'd73  : decoded = 128'b1 << 7'd73;
	7'd74  : decoded = 128'b1 << 7'd74;
	7'd75  : decoded = 128'b1 << 7'd75;
	7'd76  : decoded = 128'b1 << 7'd76;
	7'd77  : decoded = 128'b1 << 7'd77;
	7'd78  : decoded = 128'b1 << 7'd78;
	7'd79  : decoded = 128'b1 << 7'd79;
	7'd80  : decoded = 128'b1 << 7'd80;
	7'd81  : decoded = 128'b1 << 7'd81;
	7'd82  : decoded = 128'b1 << 7'd82;
	7'd83  : decoded = 128'b1 << 7'd83;
	7'd84  : decoded = 128'b1 << 7'd84;
	7'd85  : decoded = 128'b1 << 7'd85;
	7'd86  : decoded = 128'b1 << 7'd86;
	7'd87  : decoded = 128'b1 << 7'd87;
	7'd88  : decoded = 128'b1 << 7'd88;
	7'd89  : decoded = 128'b1 << 7'd89;
	7'd90  : decoded = 128'b1 << 7'd90;
	7'd91  : decoded = 128'b1 << 7'd91;
	7'd92  : decoded = 128'b1 << 7'd92;
	7'd93  : decoded = 128'b1 << 7'd93;
	7'd94  : decoded = 128'b1 << 7'd94;
	7'd95  : decoded = 128'b1 << 7'd95;
	7'd96  : decoded = 128'b1 << 7'd96;
	7'd97  : decoded = 128'b1 << 7'd97;
	7'd98  : decoded = 128'b1 << 7'd98;
	7'd99  : decoded = 128'b1 << 7'd99;
	7'd100 : decoded = 128'b1 << 7'd100;
	7'd101 : decoded = 128'b1 << 7'd101;
	7'd102 : decoded = 128'b1 << 7'd102;
	7'd103 : decoded = 128'b1 << 7'd103;
	7'd104 : decoded = 128'b1 << 7'd104;
	7'd105 : decoded = 128'b1 << 7'd105;
	7'd106 : decoded = 128'b1 << 7'd106;
	7'd107 : decoded = 128'b1 << 7'd107;
	7'd108 : decoded = 128'b1 << 7'd108;
	7'd109 : decoded = 128'b1 << 7'd109;
	7'd110 : decoded = 128'b1 << 7'd110;
	7'd111 : decoded = 128'b1 << 7'd111;
	7'd112 : decoded = 128'b1 << 7'd112;
	7'd113 : decoded = 128'b1 << 7'd113;
	7'd114 : decoded = 128'b1 << 7'd114;
	7'd115 : decoded = 128'b1 << 7'd115;
	7'd116 : decoded = 128'b1 << 7'd116;
	7'd117 : decoded = 128'b1 << 7'd117;
	7'd118 : decoded = 128'b1 << 7'd118;
	7'd119 : decoded = 128'b1 << 7'd119;
	7'd120 : decoded = 128'b1 << 7'd120;
	7'd121 : decoded = 128'b1 << 7'd121;
	7'd122 : decoded = 128'b1 << 7'd122;
	7'd123 : decoded = 128'b1 << 7'd123;
	7'd124 : decoded = 128'b1 << 7'd124;
	7'd125 : decoded = 128'b1 << 7'd125;
	7'd126 : decoded = 128'b1 << 7'd126;
	7'd127 : decoded = 128'b1 << 7'd127;
	endcase
endmodule
